magic
tech scmos
timestamp 1664280685
<< nwell >>
rect -11 24 9 30
rect -11 -7 10 24
<< polysilicon >>
rect -2 20 0 23
rect -2 -17 0 -4
rect 10 -17 12 -15
rect 22 -17 24 -15
rect 34 -17 36 -15
rect -2 -51 0 -49
rect 10 -56 12 -49
rect 22 -56 24 -49
rect 34 -56 36 -49
<< ndiffusion >>
rect -9 -29 -2 -17
rect -9 -33 -7 -29
rect -3 -33 -2 -29
rect -9 -49 -2 -33
rect 0 -49 10 -17
rect 12 -49 22 -17
rect 24 -49 34 -17
rect 36 -29 44 -17
rect 36 -33 38 -29
rect 42 -33 44 -29
rect 36 -49 44 -33
<< pdiffusion >>
rect -9 10 -2 20
rect -9 6 -7 10
rect -3 6 -2 10
rect -9 -4 -2 6
rect 0 10 8 20
rect 0 6 2 10
rect 6 6 8 10
rect 0 -4 8 6
<< metal1 >>
rect -21 32 52 36
rect -7 28 -3 32
rect -7 10 -3 24
rect 6 6 42 10
rect 38 -29 42 6
rect -7 -59 -3 -33
rect -22 -63 -7 -59
rect -3 -63 51 -59
<< ntransistor >>
rect -2 -49 0 -17
rect 10 -49 12 -17
rect 22 -49 24 -17
rect 34 -49 36 -17
<< ptransistor >>
rect -2 -4 0 20
<< polycontact >>
rect 0 -13 4 -9
rect 12 -55 16 -51
rect 24 -55 28 -51
rect 36 -55 40 -51
<< ndcontact >>
rect -7 -33 -3 -29
rect 38 -33 42 -29
<< pdcontact >>
rect -7 6 -3 10
rect 2 6 6 10
<< psubstratepcontact >>
rect -7 -63 -3 -59
<< nsubstratencontact >>
rect -7 24 -3 28
<< labels >>
rlabel polycontact 2 -11 2 -11 1 clk
rlabel metal1 40 -8 40 -8 1 out
rlabel metal1 10 -61 10 -61 1 GND
rlabel polycontact 38 -53 38 -53 1 A
rlabel polycontact 26 -53 26 -53 1 B
rlabel polycontact 14 -53 14 -53 1 C
rlabel metal1 5 34 5 34 5 VDD
<< end >>
